grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:format;

imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports silver:langutil;
imports silver:langutil:pp;

imports silver:util:treemap as tm;

