grammar determinism;

import edu:umn:cs:melt:ableC:host;

copper_mda testConcreteSyntax(ablecParser) {
  edu:umn:cs:melt:exts:ableC:halide:concretesyntax;
  edu:umn:cs:melt:exts:ableC:tensorAlgebra:concretesyntax;
}
