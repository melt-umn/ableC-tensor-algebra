grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:build;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:decls;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:format;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:indexvar;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:tensor;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:type;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:utils;
