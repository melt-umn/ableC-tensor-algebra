grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:concretesyntax;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports edu:umn:cs:melt:ableC:concretesyntax;

imports silver:langutil only ast;
