grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:env;

imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports silver:util:raw:treemap as tm;
imports silver:langutil;

global builtin::Location = builtinLoc("tensorAlgebra");
