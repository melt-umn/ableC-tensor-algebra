grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:codegen;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:syntax;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:tensors;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:type;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:env;
exports edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:expr;
