grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:indexvar;

import edu:umn:cs:melt:exts:ableC:tensorAlgebra;

abstract production indexvar
top::Decl ::= nms::[Name]
{
  local errors::[Message] =
    checkTensorHeader(head(nms).location, top.env);

  propagate substituted;
  top.pp = ppConcat([
             text("indexvar "),
             ppImplode(
               text(", "),
               map(
                 \ n::Name -> text(n.name),
                 nms)
             ),
             text(";")
           ]);

  local vars::[IndexVar] =
    map(
      \ n::Name -> indexVar(n, n.location),
      nms
    );
  
  local fwrd::Decl =
    decls(
      foldl(
        \ d::Decls v::IndexVar
        -> 
        consDecl(
          defsDecl([indexVarDef(v.variable, v)]),
          d
        )
        ,
        consDecl(
          variableDecls(
            [], 
            nilAttribute(), 
            directTypeExpr(
              indexVarType(head(nms).location)
            ),
            foldl(
              \ d::Declarators nm::Name
              -> consDeclarator(
                   declarator(nm, baseTypeExpr(), nilAttribute(), nothingInitializer()), 
                   d
                 )
              ,
              nilDeclarator(),
              nms
            )
          ),
          nilDecl()
        ),
        vars
      )
    );
  
  forwards to
  if !null(errors)
  then warnDecl(errors)
  else fwrd;
}
