grammar well_definedness;

import edu:umn:cs:melt:ableC:host;
import edu:umn:cs:melt:exts:ableC:tensorAlgebra;
