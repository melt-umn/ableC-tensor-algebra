grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:expr;

imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;
