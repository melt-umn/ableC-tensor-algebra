grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:tensor;

imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:env;
imports edu:umn:cs:melt:ableC:abstractsyntax:host;

imports edu:umn:cs:melt:exts:ableC:tensorAlgebra;

imports silver:langutil;
imports silver:langutil:pp;
