grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:expr;

