grammar edu:umn:cs:melt:exts:ableC:tensorAlgebra:abstractsyntax:decls;

imports edu:umn:cs:melt:ableC:abstractsyntax:host;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction;
imports edu:umn:cs:melt:ableC:abstractsyntax:overloadable as ovrld;
